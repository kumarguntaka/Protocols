`ifndef tb_pkg
`define tb_pkg
`include "uvm_macros.svh"
package tb_pkg;
import uvm_pkg::*;
	`include "1.transaction.sv"
	`include "2.sequence.sv"
	`include "3.driver.sv"
	`include "4.monitor.sv"
	`include "5.agent.sv"
	`include "6.scoreboard.sv"
	`include "7.environment.sv"
	`include "8.test.sv"
endpackage
`endif